library verilog;
use verilog.vl_types.all;
entity testbench_operation3 is
end testbench_operation3;
